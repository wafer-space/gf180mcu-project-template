module gf180mcu_ws_ip__id;
endmodule
